`timescale 1ns/1ns
module adder16(input[15:0] x1,x2, output[15:0] data);
    assign data = x1 + x2;
endmodule