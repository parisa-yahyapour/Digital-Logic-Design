`timescale 1ns/1ns
module multiplier16(input [15:0] x1,x2, output [15:0] result);
    assign result = x1 * x2;
endmodule